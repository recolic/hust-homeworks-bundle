/*
 * Copyright 2018-2018 Recolic Keghart <root@recolic.net>
 * Licensed under GPL 3.0
 */



