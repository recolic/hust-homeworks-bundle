
`define USE_DIVIDER
`define py