ram[0] <= 3;
ram[1] <= 1;

ram[3] <= 14;
ram[4] <= 2;

ram[6] <= 16;
ram[7] <= 4;

ram[9] <= 8'hff;
ram[10] <= 6;



ram[14] <= 6;
ram[15] <= 3;
ram[16] <= 9;
ram[17] <= 5;
